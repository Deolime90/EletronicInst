SMALL SAMPLE CIRCUIT

#REVISION: Rev: 58

.INC Pontes.MIS
V1 1 0 5 
R1 1 D  120  
R2 1 B  2400  
R3 D 0  60  
R4 B 0  1200  

* TopSpice Schematic 8.86f   Simulation Setup Commands
.DC R1 50 150 0.12
.TRAN 0.0001 0.01
.PROBE
.PRINT TRAN/ALL V(IN) D(IN) D(A) V(OUT)

.OPTION SAVEOPB
#AUTOPLOT  {V(B)-V(D)}


.END
