SMALL SAMPLE CIRCUIT

#REVISION: Rev: 97

.INC "Pontes 2.MIS"
V1 1 0 5 
R2 1 B  2400  
R3 D 0  60  
R4 B 0  1200  
X1 D 1  THERMISTOR  

* TopSpice Schematic 8.86f   Simulation Setup Commands
.DC V1 0 5 1
.STEP LIN TEMP 10 60 10
.PROBE
.PRINT TRAN/ALL V(IN) D(IN) D(A) V(OUT)

.OPTION SAVEOPB
#AUTOPLOT  {V(B)-V(D)}


.END
